`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   16:11:40 10/24/2021
// Design Name:   gray
// Module Name:   F:/sophomore/teaching assistant/ISE/P1/gray_tb.v
// Project Name:  P1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: gray
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module gray_tb;

	// Inputs
	reg Clk;
	reg Reset;
	reg En;

	// Outputs
	wire [2:0] Output;
	wire Overflow;

	// Instantiate the Unit Under Test (UUT)
	gray uut (
		.Clk(Clk), 
		.Reset(Reset), 
		.En(En), 
		.Output(Output), 
		.Overflow(Overflow)
	);
	always #5 Clk=~Clk;
	
	initial begin
		// Initialize Inputs
		Clk = 0;
		Reset = 0;
		En = 1;
		// Wait 100 ns for global reset to finish
		#105;
      Reset=1'b1;
		
		#7;	Reset=1'b0;
		
		#100	Reset=1'b1;
		
		#10	Reset=1'b0;
		// Add stimulus here

	end
      
endmodule

